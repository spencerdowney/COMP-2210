s
compiler setups
empty
      !D  "T   8
