SVe0
SVi0
SVz0
SVf0
SVj0
SVA0
SVg0
SVk0
SVB0
SVh0
SVl0
SVC0
SVp0
SVr0
SVD0
SVw0
SVy0
SVF0
SVI0
SVJ0
SVw0
SVx0
SVy0
SVF0
